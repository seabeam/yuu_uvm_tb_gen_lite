`ifndef {{ module.upper() }}_DEFINES_SVH
`define {{ module.upper() }}_DEFINES_SVH

  `ifndef {{ module.upper() }}_SETUP_TIME
  `define {{ module.upper() }}_SETUP_TIME  0
  `endif

  `ifndef {{ module.upper() }}_HOLD_TIME
  `define {{ module.upper() }}_HOLD_TIME  0
  `endif

`endif